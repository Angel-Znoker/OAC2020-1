library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
Port ( 
	dir : in STD_LOGIC_VECTOR (11 downto 0);
	data : out STD_LOGIC_VECTOR (93 downto 0));
end memory;

architecture Behavioral of memory is

begin
	process(dir)
	begin
	
		-- DATA FORMAT
		-- |    PRUEBA    |VF| Ins |                LIGA                 |
		--  P4 P3 P2 P1 P0 VF I1 I0 L11 L10 L9 L8 L7 L6 L5 L4 L3 L2 L1 L0 nCRI EB1 EB0 nWB EA1 EA0 nWA selbus UPA9 UPA8 UPA7 UPA6 UPA5 UPA4 UPA3 UPA2 UPA1 UPA0 nOEUPA nDUPA selmux nEX2 nEX1 nEX0 X2 X1 X0 EnaY nERA2 nERA1 nERA0 RA2 RA1 RA0 nEAP2 nEAP1 nEAP0 AP2 AP1 AP0 nEPC2 nEPC1 nEPC0 PC2 PC1 PC0 nCBD nAS nRW BD DINT HINT SET_IRQ SET_XIRQ B9 B8 B7 B6 B5 B4 B3 B2 B1 B0 CC CN CV CZ CI CH CX CS nHB ACCSEC

		-- Cadena por default: "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010"
		
		--if(dir=    X"000") then data <= "00000" & "0" & "00" & "000000000000" & "10010010000000000011011100001110001110001110001110000000000000000000000010";
		--elsif(dir= X"001") then data <= "00000" & "0" & "00" & "000000000000" & "00000000000000000000000000000000000000000000000000000000000000000000000000"; 
												  
												  
													-- nCRI,nWB,nWA,nOEUPA,nDUPA,nEX2,nEX1,nEX0,nERA2,nERA1,nERA0,nEAP2,nEAP1,nEAP0,nEPC1,nEPC0,nAS,nRW,nHB		
													-- Todas son negadas, por lo que están desactivadas. Las unicas banderas que están activas son
													-- nCBD y nEPC2
													-- nCRI, PC0,nAS
													-- I1, 
		if(dir=    X"000") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"001") then data <= "0000000000000000000000010010000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"002") then data <= "0000001000000000000010010010000000000011011100001110001110001110001110000000000000000000000010";

		-- LDAA #$02 Load Accumulator A
		elsif(dir= X"860") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"861") then data <= "0000000000000000000010010100000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"862") then data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000010011000000000010";
		elsif(dir= X"863") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
		elsif(dir= X"864") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

		-- LDAB #$00 Load Accumulator B
		elsif(dir= X"C60") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"C61") then data <= "0000000000000000000010100010000000000011011100001110001110001110011010000000000000000000000010";
		elsif(dir= X"C62") then data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000100101000000000010";
		elsif(dir= X"C62") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
		elsif(dir= X"C63") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

		-- ABA Add accumulator A and accumulator B
		elsif(dir= X"1B0") then data <= "0000000000000000000011111110000000000111111100001110001110001110001110000000000000000000000010";
		elsif(dir= X"1B1") then data <= "0000000000000000000010010100000000000000011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"1B2") then data <= "0111111100000000000010010010000000000010011100001110001110001110001110000000000000001111010010";
		elsif(dir= X"1B3") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

		-- JPM #$0004
		elsif(dir= X"7E0") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"7E1") then data <= "0000000000000000000010010010000000000011011100001011001110001110011011000000000000000000000010";
		elsif(dir= X"7E2") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"7E3") then data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"7E4") then data <= "0111111100000000000010010010000000000011011100001000001110001001011110000000000000000000000010";
		elsif(dir= X"7E5") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		
		-- STAA #dir
		elsif(dir= X"A70") then data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"A71") then data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
		elsif(dir= X"A72") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"A73") then data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"A74") then data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		elsif(dir= X"A75") then data <= "0000000000000000000010010110000000000011011100001110001110001110001000000000000000000000000010";
		elsif(dir= X"A76") then data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000010011000000000010";
		elsif(dir= X"A77") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
		elsif(dir= X"A78") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		
		-- GTAA #dir
		elsif(dir= X"B30") then data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"B31") then data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
		elsif(dir= X"B32") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"B33") then data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"B34") then data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		elsif(dir= X"B35") then data <= "0000000000000000000010010100000000000011011100001110001110001110001010000000000000000000000010";
		elsif(dir= X"B36") then data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000010011000000000010";
		elsif(dir= X"B37") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000010011000111000010";
		elsif(dir= X"B38") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";

		-- GTAB #dir
		elsif(dir= X"C30") then data <= "0000000000000000000010011110000100000011011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"C31") then data <= "0000000000000000000010010010000000000000011100001011001110001110001110000000000000000000000010";
		elsif(dir= X"C32") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"C33") then data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"C34") then data <= "0000000000000000000010010010000000000011011100000110001110001110000110000000000000000000000010";
		elsif(dir= X"C35") then data <= "0000000000000000000010100010000000000011011100001110001110001110001010000000000000000000000010";
		elsif(dir= X"C36") then data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000100101000000000010";
		elsif(dir= X"C37") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000100101000111000010";
		elsif(dir= X"C38") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		
		-- CBA (Acceso inherente) N,Z,V,C
		elsif(dir= X"120") then data <= "0000000000000000000011111110001010000111111100001110001110001110001110000000000000000000000011"; -- EB1,EB0,EA1,EA0,UPA7,UPA5,UPA0,selmux,ACCSEC
		elsif(dir= X"121") then data <= "0000000000000000000010010010000000000001011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"122") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000000000001111000010"; -- cc,cv,cn,cz,Prueba=15(Int), MI=11
		elsif(dir= X"123") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010"; -- Salto condicional, Prueba=24(Vale 0), es un salto forzado a la direccion x"001" y PC=Pc+1,PC0,nCBD

		-- JE #dir
		elsif(dir= X"8E0") then data <= "1001000110001110100010010010000000000011011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"8E1") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"8E2") then data <= "0000000000000000000010010010000000000011011100001011001110001110011011000000000000000000000010";
		elsif(dir= X"8E3") then data <= "0000000000000000000010010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"8E4") then data <= "0000000000000000000010010010000000000011011100001100111110001110011010000000000000000000000010";
		elsif(dir= X"8E5") then data <= "0000000000000000000010010010000000000011011100001000001110001001011110000000000000000000000010";
		elsif(dir= X"8E6") then data <= "0111111100000000000010010010000000000011011100001110001110001110001110000000000000000000000010";
		elsif(dir= X"8E7") then data <= "1100000100000000000110010010000000000011011100001110001110000110000110000000000000000000000010";
		elsif(dir= X"8E8") then data <= "0000000000000000000010010010000000000011011100001110001110001110011110000000000000000000000010";
		elsif(dir= X"8E9") then data <= "1100000110001110011010010010000000000011011100001110001110001110011110000000000000000000000010";
		
		else data <= "0000000000000000000010010010000000000011011100001110001110001110001110000000000000000000000010"; -- Default
		end if;
	end process;
end Behavioral;